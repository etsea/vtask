module task

pub struct Task {
pub:
	id int
	title string
}

pub struct TaskRepository {
	file_path string
}
